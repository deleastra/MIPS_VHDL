LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
USE ieee.numeric_std.ALL;

ENTITY instructions_memory IS
  PORT ( instruction_addr  : IN  STD_LOGIC_VECTOR(31 DOWNTO 0);
         instruction       : OUT STD_LOGIC_VECTOR(31 DOWNTO 0));
END ENTITY instructions_memory;

ARCHITECTURE dataflow OF instructions_memory IS
    TYPE mem_array IS ARRAY(31 DOWNTO 0) OF STD_LOGIC_VECTOR(31 DOWNTO 0);
	 SIGNAL instruction_mem : mem_array := (
	 "00000000000000000000000000000000", -- 0
	 "00000000000000000000000000000000",
	 "00000000000000000000000000000000",
	 "00000000000000000000000000000000",
	 "00000000000000000000000000000000",
	 "00000000000000000000000000000000",
	 "00000000000000000000000000000000",
	 "00000000000000000000000000000000",
	 "00000000000000000000000000000000",
	 "00000000000000000000000000000000",
	 "00000000000000000000000000000000", -- 10
	 "00000000000000000000000000000000",
	 "00000000000000000000000000000000",
	 "00000000000000000000000000000000",
	 "00000000000000000000000000000000",
	 "00000000000000000000000000000000",
	 "00000000000000000000000000000000",
	 "00000000000000000000000000000000",
	 "00000000000000000000000000000000",
	 "00000000000000000000000000000000",
	 "00000000000000000000000000000000", -- 20
	 "00000000000000000000000000000000",
	 "00000000000000000000000000000000",
	 "00000000000000000000000000000000",
	 "00000000000000000000000000000000",
	 "00000000000000000000000000000000",
	 "00000000000000000000000000000000",
	 "00000000000000000000000000000000",
	 "00000000000000000000000000000000",
	 "00000000000000000000000000000000",
	 "00000000000000000000000000000000",
	 "00000000000000000000000000000000"); -- 31
BEGIN
    instruction <= instruction_mem(TO_INTEGER(UNSIGNED(instruction_addr)));
END dataflow;